// Code your testbench here
// or browse Examples
module tb;
  initial
    begin
    	$display("HELLO WORLD,I m verilog");
    end
endmodule
